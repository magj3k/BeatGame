BZh91AY&SY��Es s_�Px����߰����POt���*(H�H�B��LB2jyd�51C��)�mR�� ���  4Ч��zP��z�     9�&L�0�&&��!�0# �54'��6�i0�j  L��@Cs �������	?����(6X�h d5�d��젒/E�]M� �����P�M<3؊���OM&tU�k��ƹ ��%Cybb���˶~ǫaݍ	*o�_���uC6B�`��En.���(GЁ�0Ɇ����f��g\��E�eѻ9���H!���fm&��p�H�� EFw/��(g8���-c$�a�:C�8ʰ�СR�qk�A2�3��ZPtT��{*KC	5��T�H��A��Q�!=bBJ��f��Z�,ڑZ�m*6�D�c���3		9D�@( �ݜ���y*M
.J�e�ԗ5A��hH�2@4�B�(9�U2�npvPe�*�t fQn.�6���D��'�O]�UR�>R~c[v8w��Œ�U��g�/J"&��+���w.����m�iZ}�����n���@t,��c��7'�Q�8u�.��T�8���E�!2���:�D�'�TY��~�N�r]u��!��S&.a�^\��:1�x��i)pm���YwG�C2;yL��{��ƃ�����o�~��FCˬ���)�|�Ӆ00 {��_Q�N��+1!|R ��q�^jR]�P�36�������NM��4*��ǅ0����H�ss�"b���|R֊��h`Yk*Ł(�Je�W	�(��{��I�������@0X)��c-%�\y
�@�P~z�܂�-AI(��R;�\g̷֜Y�9q\N܃h,��΃Q_:�T l�I�w�o�!%�%iE�Vȋ�*�7��Q�U�i��έ!l�{x�{��P���U�����Ŭ��d#IP�}��>��C�PwF7؆����)�n�qcu�Ƅ3.%��ƓC%���S]�w$S�		)�W0