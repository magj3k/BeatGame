BZh91AY&SYr�{� �߀Px����߰����P�r��1@$�4�OI�����P i� �@jz$f�I4�� ��   M4P�� �6�� di�A��bdɣ	�bi�L#0	&�M�E1'���=L���OS�M.�!�DJ����_&C!��	O��v�<Xb^ ��&�;�!Z4����9 PZ�~�ݶl��4,���@����J�W�@�a��p����uk��!"�����a�Lѫ�-�a$ R�	$
��w�|c��d�^�U�Qd��Z��"[��s�L�gY���VX�J�8�p���;�	&N�8@92�`m�3=�Q5JX"��Dā�YPZ)J:D�K
�EK.l�I�ւ�tp�r,Z�A�MĒ@0  Aѵy�]�? y
6��G�B*@�M(RZ�C���d�m���ɦ@J-���PԚ����$aS���t�v��
nb��оg)�Ņt��ۇ*�~�����|Z�DSrYǸ���_��)��1���d�\@��83)���)�QRp�Gq�\��g"��8(�B�f�- z,D�F�.:Gu} ��檪��pԧf.P�
.�)���pg(Ф��RM]d>�؂P����D�� �
kĠI���خd6k��Ȣ�TK�J;'ϭ0`�!~=�~j�U�q#&$���ii���_YC1���r�\b+0l{׎
����0��-0i �I�ys�Y5�����в(Ũ�/��� �\�QD%�(
}��$�(�c�dLV*U3�er*�j��A)�o�uf!����H[o-!����~���14�o�>p��g�y��Ȭ��oLkoN�ES$�D�櫱6Qn��8Lv��*3V���m�x�TTJ�2V�0
Y�"�cZ@�E��� �l�HF=Q��i�P��N���
���jr���2�R�]2�Y���rE8P�r�{�