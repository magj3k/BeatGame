BZh91AY&SYqp� �_�Px����߰����P��n��6�A�E )�T�Bm��j4��2$=M=OP��j~T��F�    DD�4��@4�'���Q� �=&C�bdɣ	�bi�L#0	$�4`T��=F�z��  h�U �Q%`G��(%;�>���X� L��Q�($`4���5����5���6eqӵ,�ܟ��I|(��1��Qv��u���f1�aiN�LK�$J�a{t$�A��H�<��]đ��y9_��:�ݩrh�V�}��HL��Q��OL�04i`Yl���	�j؈�9���V��X�Ёa�Q X�d����c��D	�$9�ݶ�������61���m�hPAùʷB44 �4(��f_������h,˥���F�^PR�K�!�kՋ�hM���!����g�)�5^�v���>�c��I<=䄤���dV���h� ��W�|�� [�i�3"��Fk�WOQ�o������	@9����!8l�q���ݡx�҅/�PrF�D�'C.b�k�������7��	Ќ��[3���a�2��}z]�rl!"`���֨�!��tI�8w�GP���&��U"=P��x��ԞLI'
�wK���D�"��&\��?b�A!����ЃF�Ӑ��4Q'�H�[�W�K:�=83�|�����0�Di"�Z��Bb��o{��%Q�/&��&��Ƽ�| �	��9�z�D���|?|P�Jnfc-%�*�BPQoېCi�@�Gv�`�t�Ĥ<��@\(��u����0d m�ػ�U&�pL2ӣPX�Du�7��(�14@�����j���jL_�~�T�'Y�ր�B����
T����&V�F��T��7>�	!�l���C� eAۨ�uA����\3�m~�T�w�Q�KYi���"�(H8�� 