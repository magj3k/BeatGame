BZh91AY&SY�ֵ �_�Px����߰����P�t]p�Ѩ$�4&&)��OR`@�F "��OJ   hh�  ��5MOj&��j0LF�a 4ɑ��9�&L�0�&&��!�0# �Ade57�S&�=� ��� = " 
bJ�G�"P�x}� �6ؗp&A��8d��ƑC֠�����sFYh�k�I�O����m���B6��Äq���ȉ3�ۉ���X>|�9}�C)�W�qBJVQ��H�=}tf�L�	�1���o�GW"��qj*��D�1���P��Ж�R@b�ɰ_Bz�,Zj�mb+:�i��8�k� P�� �12H�
&��DBZ�A��6��һ�1��f3p��"�䪃I'g�r=��	31�S.��\LIc��JT�!��BK��d%��3��ac&�s�mn�<���WF�t*d5v?չ����]�	4�˕������P)j�̿`���h�J�!iW_f+���(�][/�}Tgn"���ę�x�|��]�4!K�ur^VC8��j�I�5����|���rQE5��lʥV0dk}S�jH�Ѥip5
)�!6A��xD2#���\V���c�^*��I�WƼ�fj��ɨ�8*Imʏ	1�00'Dr��I�;��+�#�K�E�.�+/Q(�H�3&_y<���Vfǭp̦9�:���Z�" �w�0���mײ� l�d�96,�Ql�e�yc"(���D	&NDo/�l�jEb�"^�fX���Dłu�:q�� ^�\ą���<w�HtXj�r����e���|��@΍���*�!^l#�"	�q�b �D��"�*jE���ipLy�u�Wm��)�Pa��R��H?�`
VZ� C%�Z��0&�M!=c�}���"����7X�*���l�e3�F�_�d*Y��	��Œ���(�?�]��BC��Z�