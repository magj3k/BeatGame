BZh91AY&SY�A�j �_�Px����߰����P�wn����*�:�I"���&��D�2!�  h	B&L�I���� @ � �4z��4�  444�ɓF�� �0F`( O�Jzi�M��T� b��E� {@D ĕ ��P0$%�����6%� ��8l��ƑCmA�BkS^�$$�lC^�(Eơ����L�B�5��ߎ��]���TXP{FLHZ1aDyls��U$�A��-gd��L�c�\|h�D�8ֶE%�;��m:�.�d��3��I�DC"�j�j�F������Ib
����TZ�����G�礦麐��%r���QY�RO���U�W��l��VU�/lccn��`Р@���Y��C�"D����B��j�7C�	���f�D�dB� TptЛ�˴v$��3X��5p�W��Ù,y���kʸ0�v|����KCei��X��U�PUJ��'�P����*˘�wcԊ��e_����癆�f�(���ڻFmB�`��܏�5f�-!�&{fخ�|u��>
R�+|��iY����6��&091 
.B�j�M�y��Z�B�A;(&uEx��I8M�����4ĂxH?��vZ�R``NEec����&䚔o�+�`��=�l+/JE>�f#.�,����P(�{c�k��4-G
`{�N]d�Yw��aa�F��UAV���dش�Eҕ��	��L�ĂY?��L���c�ǐ��E����Hrr��p���>�YG�4�`��({��@X���h��`��9�9�URB|i&5���
��D���#*jE�D�Qd`�ؒ�/_��D��3.��,����
u �fZ��/&U�HO!��($M�H4�DjCjR��	��#b��_��/��	|)3�l(*��]��BB)ɨ