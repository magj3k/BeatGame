BZh91AY&SY"�? �_�Px����߰����P�wn��8U(P�DИ��ވS�)�����i�zP��2�~BM��4      �J�ڀ f�     昙2h�`��` ���D� ML��L�i�Ȟ�# 4���4�@�!�B� �H��2<R~�8�;�Ļ��w��}j�ib�J��6.Y���a.��JP�y�SNER�r_�	U�!��b9�B|D>AI�{ZB�� Q���
���<b�͓D�S}"��y��É&q&0�y����-�W�#����s[3@�h{ͣ<���K%����YRX2����A��/k,%U�x�Ȋ��lݮ5�J����LR����a�6���d�B2�	4_J�hj����c�B@ �ۅ�G]��[��j"d��T��S ���
1�Jb�j)T%���J`�>�)n��<�y���<2�o�������HI}��·���1]�y_d�#�x�q�%z�u�m>�]̼<��<K򜓃j��ۈ�Oɜ��G���3��^�.���� �3��1��*�����wvu#�ֻ��<ʷ�����|��X�:|$$R�XĲ_��P����(f`��IƳz��#�@�]�ٝ�n���u�G����$�r��H�j�/b�!���Θ+����eGʥݤ�#5o?bv�n���}�+�ɡ0=����[2D��v���VA`4�d�n%���5V��'���"Ĥ.� P���(S%@ǌ?TT��g�2��jǐ�������lq�K�x���9���Y8|�ۚ�q���x�ƂH8�;�
���#�c[���l
�E�W^�l�o�P&<~xڥ��6�u+�bn�R��$*Sj%7��v��B6�\�~-v%;��}U[b�qЃ�9	T�'"��9s�K2�P��T�\X4��.�p� 4E�~