BZh91AY&SY�k� u_�Px����߰����P�v���	$ ��������)��� �ڟ�h�2?Ri��&�&	��0`��4��
��bh�M   9�&L�0�&&��!�0# �#D&I���B��jz�1���=H�I�D���W`�h�A(~�y2`K��k�ʮ�PF#H���`L5+��~��rL\ցI?��i�N��y�0�~�K�u?>Y�����HS��"5T-F��3���BS6ƨH�o��vsƘ�ev4U�\pY23�"s����c�,�VL����d2MHH$e��$�|�����SI�B,I����n-�QKP�[l�� ̶f�̖Tש���	�U
j1�A�	�Ӯ]}��vXy��w7��R����	}�3�� 3d�I�t�鄞S�N4�Yh�`���2��Z&ƨ�F��Z�,�Q��iݶ3s'�!��4ָ�kz4SG<dT�������i��nշy����j'���?I�87��e�xpL�<z9�KzWx��P�#Q�9:�0H�,ag��U�W~��_�����Y�j��!��0�&��y��H#�*&��d?O��P�lG��P�Łq:JJ��[��L���v#�)L!ʡ��q�f�~*�#͚0-�0m����fjqU/�I�f|�/�<28������J4��Z`{��B.��x�Z���W��+�6�K�,[J#:�-�����#� P���(S&<a��n[�,ϔe�Z!�䂅P�{��.�>r�㙉<��v�ݑ����m�f����	 ���4�5H�jSΑ	�r���-R�z0���$EY�	���8)f��?,����`�)!R�L�H�b�DA75�f2�����	�~��%<h���>=y�F/ì�ԝP�ݥ˞��e�X���6�X02��.�p�!T4�H