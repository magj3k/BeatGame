BZh91AY&SYgi �_�Px����߰����P�wn�;����	B�&�`i'���@SMA�M ���'����&    	S�J=�FM4ѧ�A�@� ѐ0昙2h�`��` ���D�	����C$ɦ�� 4��K�{�� �������|�	��F%����Y7�1
ѤT���0(�%v�EM�
�rX�q�B�?��I�<Nk�SfeP�|�_bs2���
dŀt� �1`�R����I ����
���U��� Ƙ�m�L�[���P���d�XД��
t�n:�D4J\$T6,�H�����I��mcz���pE�ÔqtC�L)3T.+8
�"��LZ��MQ�b��ž�/���B��,�:��HIn$� Ͼ���_�6�D6�ۜ&�#a�l�r���D@�<M2�U@CTj�y�Bl/fȌ�����Iɮ�?:^q��U̴��5���sғ�f��9 "�Ri���
Qq�ݎb)@5%5O�����N�YW�T�?���W�/Y�"�kN"H�4��]�7�����9�B�f,YC�����`�߼�y�X		�9�)�4��]���<�n�&��B�E$��FC���dG���e-`V �[���c�YA�ۜl�ç9E � ��,�hu�"��3�O�ɿfX����@{���ZfR*�&i�lV���0+0lz��
����L%+L�!b��s	�?�XQZ�h�g(ŴI�wf)�a:BLL%��H	�Q@�d?�L
U3�er*�j�����0�9O^���,@:�=Dū)q<�o�5�Ta1���d9���PɌ��F�p���נ0H�d�dL�5]�����E䁤�01�L�r0��鴨�R�7{L+��b� �,����A���v��
j>(��A���!��eA��)R���sD.����*���q���0h.�g�]��BA�M�h